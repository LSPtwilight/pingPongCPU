
//`include "defines.v"

`define DivIdle     2'b00
`define DivByZero   2'b01
`define DivOn       2'b10
`define DivEnd      2'b11
`define ZeroWord    32'd0

module div(
	input clk, resetn,
	
	input 	[31:0] 	    opdata1_i,
	input 	[31:0] 	    opdata2_i,
	input 				signed_div_i,
	input 				start_i,
	input 				annul_i,	// cancel division
	
	output reg 	[63:0]  result_o,
	output reg 			ready_o
);

	reg 	[64:0] 	dividend;
	wire 	[32:0] 	div_temp;
	reg 	[31:0] 	divisor;
	reg 	[5:0] 	cnt;
	reg 	[1:0] 	state;

	reg     sign_1;
	reg     sign_2;

	assign div_temp = {1'b0, dividend[63:32]} - {1'b0, divisor};

	always @ (posedge clk) begin
		if (!resetn) begin
			state 	<= `DivIdle;
			ready_o <= 1'b0;
			result_o <= {`ZeroWord,`ZeroWord};
		end else begin
		    case (state)
		  	`DivIdle: begin               //DivIdle
		  		if (start_i == 1'b1 && annul_i == 1'b0) begin
		  			if (opdata2_i == `ZeroWord) begin
		  				state <= `DivByZero;
		  			end else begin
		  				state <= `DivOn;
		  				cnt <= 6'b000000;
		  				dividend[63:33] <= 31'b0;
		  				dividend[0] <= 1'b0;
						sign_1 <= opdata1_i[31];
						sign_2 <= opdata2_i[31];
		  				if (signed_div_i == 1'b1 && opdata1_i[31] == 1'b1 ) begin
		  					dividend[32:1] <= ~opdata1_i + 1;
		  				end else begin
		  					dividend[32:1] <= opdata1_i;
		  				end
		  				if (signed_div_i == 1'b1 && opdata2_i[31] == 1'b1 ) begin
		  					divisor <= ~opdata2_i + 1;
		  				end else begin
		  					divisor <= opdata2_i;
		  				end
                     end
                end else begin
				     ready_o <= 1'b0;
					 result_o <= {`ZeroWord,`ZeroWord};
				end          	
		  	end
		  	`DivByZero:	begin               //DivByZero
         	    dividend <= {`ZeroWord,`ZeroWord};
                state <= `DivEnd;		 		
		  	end
		  	`DivOn:	begin               //DivOn
		  		if (annul_i == 1'b0) begin
		  			if (cnt != 6'b100000) begin 	// cnt reach 32
                        if (div_temp[32] == 1'b1) begin 	// 商这一位取0
                            dividend <= {dividend[63:0] , 1'b0};	// 最后跟着的一位就是商
                        end else begin
                            dividend <= {div_temp[31:0] , dividend[31:0] , 1'b1};
                        end
                    	cnt <= cnt + 1;
                    end else begin
                        if ((signed_div_i == 1'b1) && ((/*opdata1_i[31] ^ opdata2_i[31]*/sign_1 ^ sign_2) == 1'b1)) begin
                            dividend[31:0] <= (~dividend[31:0] + 1);
                        end
                        if ((signed_div_i == 1'b1) && ((/*opdata1_i[31]*/sign_1 ^ dividend[64]) == 1'b1)) begin              
                            dividend[64:33] <= (~dividend[64:33] + 1);
                        end
                    	state <= `DivEnd;
                    	cnt <= 6'b000000;
                	end
		    	end else begin
		  			state <= `DivIdle;
		  		end	
		  	end
		  	`DivEnd: begin               //DivEnd
        		result_o 	<= {dividend[64:33], dividend[31:0]};  	// 高32为余数，低32为商
          		ready_o 	<= 1'b1;
          		if (start_i == 1'b0) begin
          			state 	<= `DivIdle;
					ready_o <= 1'b0;
					result_o <= {`ZeroWord,`ZeroWord};       	
          		end		  	
		  	end
		  endcase
		end
	end
endmodule
